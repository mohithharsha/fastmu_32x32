// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_proj_example
 *
 * This is an example of a (trivially simple) user project,
 * showing how the user project can connect to the logic
 * analyzer, the wishbone bus, and the I/O pads.
 *
 * This project generates an integer count, which is output
 * on the user area GPIO pads (digital output only).  The
 * wishbone connection allows the project to be controlled
 * (start and stop) from the management SoC program.
 *
 * See the testbenches in directory "mprj_counter" for the
 * example programs that drive this user project.  The three
 * testbenches are "io_ports", "la_test1", and "la_test2".
 *
 *-------------------------------------------------------------
 */

module user_proj_example #(
    parameter BITS = 32
)(
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // IRQ
    output [2:0] irq
);
    wire clk;
    wire rst;

    wire [`MPRJ_IO_PADS-1:0] io_in;
    wire [`MPRJ_IO_PADS-1:0] io_out;
    wire [`MPRJ_IO_PADS-1:0] io_oeb;

    wire [31:0] rdata; 
    wire [31:0] wdata;
    wire [BITS-1:0] count;

    wire valid;
    wire [3:0] wstrb;
    wire [31:0] la_write;

    // WB MI A
    assign valid = wbs_cyc_i && wbs_stb_i; 
    assign wstrb = wbs_sel_i & {4{wbs_we_i}};
    assign wbs_dat_o = rdata;
    assign wdata = wbs_dat_i;

    // IO
    assign io_out = count;
    assign io_oeb = {(`MPRJ_IO_PADS-1){rst}};

    // IRQ
    assign irq = 3'b000;	// Unused

    // LA
    assign la_data_out = {{(127-BITS){1'b0}}, count};
    // Assuming LA probes [63:32] are for controlling the count register  
    assign la_write = ~la_oenb[63:32] & ~{BITS{valid}};
    // Assuming LA probes [65:64] are for controlling the count clk & reset  
    assign clk = (~la_oenb[64]) ? la_data_in[64]: wb_clk_i;
    assign rst = (~la_oenb[65]) ? la_data_in[65]: wb_rst_i;

fastmul_32x32 dut(a,b,y);

endmodule


module fastmul_32x32(a,b,y);
input [31:0]a,b;
  output [63:0]y;
  wire[1023:0]p;
  wire [180:12]s,c; 
wire[111:0]s1,c1,Cout;
wire [38:0]o0,o1,o2,o3;
wire [7:0]O0,O1,O2,O3,O4;

mul_16x16 u35(a[15:0],b[15:0],p[255:0]);
mul_16x16 u36(a[31:16],b[15:0],p[511:256]);
mul_16x16 u37(a[15:0],b[31:16],p[767:512]);
mul_16x16 u38(a[31:16],b[31:16],p[1023:768]);

//first stage
//4
ha u39(p[4],p[35],s[12],c[12]);
//5
counter53 u40(p[5],p[36],p[67],p[98],c[12],s1[0],c1[0],Cout[0]);
//6
counter53 u41(p[6],p[37],p[68],p[99],c1[0],s1[1],c1[1],Cout[1]);
//7
counter53 u42(p[7],p[38],p[69],p[100],Cout[0],s1[2],c1[2],Cout[2]);
fa u43(p[131],p[162],c1[1],s[13],c[13]);
//8
counter53 u44(p[8],p[39],p[70],p[101],Cout[1],s1[3],c1[3],Cout[3]);
counter53 u45(c1[2],c[13],p[132],p[163],p[194],s1[4],c1[4],Cout[4]);
//9
counter53 u46(p[9],p[40],p[71],p[102],Cout[2],s1[5],c1[5],Cout[5]);
counter53 u47(c1[3],c1[4],p[133],p[164],p[195],s1[6],c1[6],Cout[6]);
//10
counter53 u48(p[10],p[41],p[72],p[103],Cout[3],s1[7],c1[7],Cout[7]);
counter53 u49(Cout[4],c1[5],c1[6],p[134],p[165],s1[8],c1[8],Cout[8]);
ha u50(p[196],p[227],s[14],c[14]);
//11
counter53 u51(p[11],p[42],p[73],p[104],Cout[5],s1[9],c1[9],Cout[9]);
counter53 u52(Cout[6],c1[7],c1[8],c[14],p[135],s1[10],c1[10],Cout[10]);
fa u53(p[166],p[197],p[228],s[15],c[15]);
//12
counter154 u54(p[12],p[43],p[74],p[105],p[136],p[167],p[198],p[229],p[260],p[291],p[322],p[353],p[384],Cout[7],Cout[8],o0[0],o1[0],o2[0],o3[0]);
//13
counter154 u55(p[13],p[44],p[75],p[106],p[137],p[168],p[199],p[230],p[261],p[292],p[323],p[354],p[385],p[416],o1[0],o0[1],o1[1],o2[1],o3[1]);
//14
counter154 u56(p[14],p[45],p[76],p[107],p[138],p[169],p[200],p[231],p[262],p[293],p[324],p[355],p[386],p[417],p[448],o0[2],o1[2],o2[2],o3[2]);
//15
counter154 u57(p[15],p[46],p[77],p[108],p[139],p[170],p[201],p[232],p[263],p[294],p[325],p[356],p[387],p[418],p[449],o0[3],o1[3],o2[3],o3[3]);
ha u58(O3[0],p[480],s[16],c[16]);
//16
counter154 u59(p[16],p[47],p[78],p[109],p[140],p[171],p[202],p[233],p[264],p[295],p[326],p[357],p[388],p[419],p[450],o0[4],o1[4],o2[4],o3[4]);
fa u60(O3[1],p[481],p[512],s[17],c[17]);
//17
counter154 u61(p[17],p[48],p[79],p[110],p[141],p[172],p[203],p[234],p[265],p[296],p[327],p[358],p[389],p[420],p[451],o0[5],o1[5],o2[5],o3[5]);
fa u62(p[482],p[513],p[544],s[18],c[18]);
//18
counter154 u63(p[18],p[49],p[80],p[111],p[142],p[173],p[204],p[235],p[266],p[297],p[328],p[359],p[390],p[421],p[452],o0[6],o1[6],o2[6],o3[6]);
counter53 u64(p[483],p[514],p[545],p[576],o3[3],s1[11],c1[11],Cout[11]);
//19
counter154 u65(p[19],p[50],p[81],p[112],p[143],p[174],p[205],p[236],p[267],p[298],p[329],p[360],p[391],p[422],p[453],o0[7],o1[7],o2[7],o3[7]);
counter53 u66(p[484],p[515],p[546],p[577],p[608],s1[12],c1[12],Cout[12]);
//20
counter154 u67(p[20],p[51],p[82],p[113],p[144],p[175],p[206],p[237],p[268],p[299],p[330],p[361],p[392],p[423],p[454],o0[8],o1[8],o2[8],o3[8]);
counter53 u68(p[485],p[516],p[547],p[578],p[609],s1[13],c1[13],Cout[13]);
fa u69(p[640],o3[5],o2[6],s[19],c[19]);
//21
counter154 u70(p[21],p[52],p[83],p[114],p[145],p[176],p[207],p[238],p[269],p[300],p[331],p[362],p[393],p[424],p[455],o0[9],o1[9],o2[9],o3[9]);
counter53 u71(p[486],p[517],p[548],p[579],p[610],s1[14],c1[14],Cout[14]);
fa u72(p[641],p[672],o3[6],s[20],c[20]);
//22
counter154 u73(p[22],p[53],p[84],p[115],p[146],p[177],p[208],p[239],p[270],p[301],p[332],p[363],p[394],p[425],p[456],o0[10],o1[10],o2[10],o3[10]);
counter53 u74(p[487],p[518],p[549],p[580],p[611],s1[15],c1[15],Cout[15]);
fa u75(p[642],p[673],p[704],s[21],c[21]);
//23
counter154 u76(p[23],p[54],p[85],p[116],p[147],p[178],p[209],p[240],p[271],p[302],p[333],p[364],p[395],p[426],p[457],o0[11],o1[11],o2[11],o3[11]);
counter53 u77(p[488],p[519],p[550],p[581],p[612],s1[16],c1[16],Cout[16]);
fa u78(p[643],p[674],p[705],s[22],c[22]);
//24
counter154 u79(p[24],p[55],p[86],p[117],p[148],p[179],p[210],p[241],p[272],p[303],p[334],p[365],p[396],p[427],p[458],o0[12],o1[12],o2[12],o3[12]);
counter53 u80(p[489],p[520],p[551],p[582],p[613],s1[17],c1[17],Cout[17]);
fa u81(p[644],p[675],p[706],s[23],c[23]);
//25
counter154 u82(p[25],p[56],p[87],p[118],p[149],p[180],p[211],p[242],p[273],p[304],p[335],p[366],p[397],p[428],p[459],o0[13],o1[13],o2[13],o3[13]);
counter53 u83(p[490],p[521],p[552],p[583],p[614],s1[18],c1[18],Cout[18]);
fa u84(p[645],p[676],p[707],s[24],c[24]);
//26
counter154 u85(p[26],p[57],p[88],p[119],p[150],p[181],p[212],p[243],p[274],p[305],p[336],p[367],p[398],p[429],p[460],o0[14],o1[14],o2[14],o3[14]);
counter53 u86(p[491],p[522],p[553],p[584],p[615],s1[19],c1[19],Cout[19]);
fa u87(p[646],p[677],p[708],s[25],c[25]);
//27
counter315 u88(p[27],p[58],p[89],p[120],p[151],p[182],p[213],p[244],p[275],p[306],p[337],p[368],p[399],p[430],p[461],p[492],p[523],p[554],p[585],p[616],p[647],p[678],p[709],p[740],p[771],p[802],p[833],p[864],o3[12],o2[13],Cout[18],O0[0],O1[0],O2[0],O3[0],O4[0]);
ha u89(o1[14],c1[19],s[26],c[26]);
//28
counter315 u90(p[28],p[59],p[90],p[121],p[152],p[183],p[214],p[245],p[276],p[307],p[338],p[369],p[400],p[431],p[462],p[493],p[524],p[555],p[586],p[617],p[648],p[679],p[710],p[741],p[772],p[803],p[834],p[865],p[896],O1[0],c[26],O0[1],O1[1],O2[1],O3[1],O4[1]);

//29
counter315 u91(p[29],p[60],p[91],p[122],p[153],p[184],p[215],p[246],p[277],p[308],p[339],p[370],p[401],p[432],p[463],p[494],p[525],p[556],p[587],p[618],p[649],p[680],p[711],p[742],p[773],p[804],p[835],p[866],p[897],p[928],O2[0],O0[2],O1[2],O2[2],O3[2],O4[2]);
//30
counter315 u92(p[30],p[61],p[92],p[123],p[154],p[185],p[216],p[247],p[278],p[309],p[340],p[371],p[402],p[433],p[464],p[495],p[526],p[557],p[588],p[619],p[650],p[681],p[712],p[743],p[774],p[805],p[836],p[867],p[898],p[929],p[960],O0[3],O1[3],O2[3],O3[3],O4[3]);
//31
counter315 u93(p[31],p[62],p[93],p[124],p[155],p[186],p[217],p[248],p[279],p[310],p[341],p[372],p[403],p[434],p[465],p[496],p[527],p[558],p[589],p[620],p[651],p[682],p[713],p[744],p[775],p[806],p[837],p[868],p[899],p[930],p[961],O0[4],O1[4],O2[4],O3[4],O4[4]);
//32
counter315 u94(p[63],p[94],p[125],p[156],p[187],p[218],p[249],p[280],p[311],p[342],p[373],p[404],p[435],p[466],p[497],p[528],p[559],p[590],p[621],p[652],p[683],p[714],p[745],p[776],p[807],p[838],p[869],p[900],p[931],p[962],p[993],O0[5],O1[5],O2[5],O3[5],O4[5]);
//33- 30 e
counter315 u95(p[95],p[126],p[157],p[188],p[219],p[250],p[281],p[312],p[343],p[374],p[405],p[436],p[467],p[498],p[529],p[560],p[591],p[622],p[653],p[684],p[715],p[746],p[777],p[808],p[839],p[870],p[901],p[932],p[963],p[994],O4[2],O0[6],O1[6],O2[6],O3[6],O4[6]);
//34 -29 e
counter315 u96(p[127],p[158],p[189],p[220],p[251],p[282],p[313],p[344],p[375],p[406],p[437],p[468],p[499],p[530],p[561],p[592],p[623],p[654],p[685],p[716],p[747],p[778],p[809],p[840],p[871],p[902],p[933],p[964],p[995],O4[3],O3[4],O0[7],O1[7],O2[7],O3[7],O4[7]);
//35 -28 e
counter154 u97(p[159],p[190],p[221],p[252],p[283],p[314],p[345],p[376],p[407],p[438],p[469],p[500],p[531],p[562],p[593],o0[15],o1[15],o2[15],o3[15]);
counter154 u98(p[624],p[655],p[686],p[717],p[748],p[779],p[810],p[841],p[872],p[903],p[934],p[965],p[996],O4[4],O3[5],o0[16],o1[16],o2[16],o3[16]);
//36 -27 e
counter154 u99(p[191],p[222],p[253],p[284],p[315],p[346],p[377],p[408],p[439],p[470],p[501],p[532],p[563],p[594],p[625],o0[17],o1[17],o2[17],o3[17]);
counter154 u100(p[656],p[687],p[718],p[749],p[780],p[811],p[842],p[873],p[904],p[935],p[966],p[997],O4[5],O3[6],O2[7],o0[18],o1[18],o2[18],o3[18]);
//37 -26 e
counter154 u101(p[223],p[254],p[285],p[316],p[347],p[378],p[409],p[440],p[471],p[502],p[533],p[564],p[595],p[626],p[657],o0[19],o1[19],o2[19],o3[19]);
counter154 u102(p[688],p[719],p[750],p[781],p[812],p[843],p[874],p[905],p[936],p[967],p[998],O4[6],O3[7],o2[15],o2[16],o0[20],o1[20],o2[20],o3[20]);
//38 -25 e
counter154 u103(p[255],p[286],p[317],p[348],p[379],p[410],p[441],p[472],p[503],p[534],p[565],p[596],p[627],p[658],p[689],o0[21],o1[21],o2[21],o3[21]);
counter154 u104(p[720],p[751],p[782],p[813],p[844],p[875],p[906],p[937],p[968],p[999],O4[7],o3[15],o3[16],o2[17],o2[18],o0[22],o1[22],o2[22],o3[22]);
//39 - 24 e
counter154 u105(p[287],p[318],p[349],p[380],p[411],p[442],p[473],p[504],p[535],p[566],p[597],p[628],p[659],p[690],p[721],o0[23],o1[23],o2[23],o3[23]);
counter154 u106(p[752],p[783],p[814],p[845],p[876],p[907],p[938],p[969],p[1000],o3[17],o3[18],o2[19],o2[20],o1[21],o1[22],o0[24],o1[24],o2[24],o3[24]);
//40 -23 e
counter154 u107(p[319],p[350],p[381],p[412],p[443],p[474],p[505],p[536],p[567],p[598],p[629],p[660],p[691],p[722],p[753],o0[25],o1[25],o2[25],o3[25]);
counter53 u108(p[784],p[815],p[846],p[877],p[908],s1[20],c1[20],Cout[20]);
counter53 u109(p[939],p[970],p[1001],o3[19],o3[20],s1[21],c1[21],Cout[21]);
//41 -22 e
counter154 u110(p[351],p[382],p[413],p[444],p[475],p[506],p[537],p[568],p[599],p[630],p[661],p[692],p[723],p[754],p[785],o0[26],o1[26],o2[26],o3[26]);
counter53 u111(p[816],p[847],p[878],p[909],p[940],s1[22],c1[22],Cout[22]);
  counter53 u112(p[971],p[1002],o3[21],o3[22],o2[23],s1[23],c1[23],Cout[23]);
//42 -21 e
  counter154 u113(p[383],p[414],p[445],p[476],p[507],p[538],p[569],p[600],p[631],p[662],p[693],p[724],p[755],p[786],p[817],o0[27],o1[27],o2[27],o3[27]);
  counter53 u114(p[848],p[879],p[910],p[941],p[972],s1[24],c1[24],Cout[24]);
  counter53 u115(p[1003],o3[23],o3[24],o2[25],Cout[20],s1[25],c1[25],Cout[25]);
//43 -20 e
  counter154 u116(p[415],p[446],p[477],p[508],p[539],p[570],p[601],p[632],p[663],p[694],p[725],p[756],p[787],p[818],p[849],o0[28],o1[28],o2[28],o3[28]);
  counter53 u117(p[880],p[911],p[942],p[973],p[1004],s1[26],c1[26],Cout[26]);
  counter53 u118(o3[25],o2[26],Cout[22],Cout[23],o1[27],s1[27],c1[27],Cout[27]);

  
//44 -19 e
counter154 u119(p[447],p[478],p[509],p[540],p[571],p[602],p[633],p[664],p[695],p[726],p[757],p[788],p[819],p[850],p[881],o0[29],o1[29],o2[29],o3[29]);
counter53 u120(p[912],p[943],p[974],p[1005],o3[26],s1[28],c1[28],Cout[28]);
counter53 u121(o2[27],Cout[24],Cout[25],o1[28],c1[26],s1[29],c1[29],Cout[29]);
//45 - 18 e
counter154 u122(p[479],p[510],p[541],p[572],p[603],p[634],p[665],p[696],p[727],p[758],p[789],p[820],p[851],p[882],p[913],o0[30],o1[30],o2[30],o3[30]);
counter53 u123(p[944],p[975],p[1006],o3[27],o2[28],s1[30],c1[30],Cout[30]);
counter53 u124(Cout[26],Cout[27],o1[29],c1[28],c1[29],s1[31],c1[31],Cout[31]);
//46 - 17 e
counter154 u125(p[511],p[542],p[573],p[604],p[635],p[666],p[697],p[728],p[759],p[790],p[821],p[852],p[883],p[914],p[945],o0[31],o1[31],o2[31],o3[31]);
counter53 u126(p[976],p[1007],o3[28],o2[29],Cout[28],s1[32],c1[32],Cout[32]);
fa u127(Cout[29],o1[30],c1[30],s[26],c[26]);
//47 - 16 e
counter154 u128(p[543],p[574],p[605],p[636],p[667],p[698],p[729],p[760],p[791],p[822],p[853],p[884],p[915],p[946],p[977],o0[32],o1[32],o2[32],o3[32]);
counter53 u129(p[1008],o3[29],o2[30],Cout[30],Cout[31],s1[33],c1[33],Cout[33]);
ha u130(o1[31],c1[32],s[27],c[27]);
//48 - 15 e
counter154 u131(p[575],p[606],p[637],p[668],p[699],p[730],p[761],p[792],p[823],p[854],p[885],p[916],p[947],p[978],p[1009],o0[33],o1[33],o2[33],o3[33]);
counter53 u132(o3[30],o2[31],Cout[32],o1[32],c1[33],s1[34],c1[34],Cout[34]);
//49 - 14 e
counter154 u133(p[607],p[638],p[669],p[700],p[731],p[762],p[793],p[824],p[855],p[886],p[917],p[948],p[979],p[1010],o3[31],o0[34],o1[34],o2[34],o3[34]);
fa u134(o2[32],Cout[33],o1[33],s[28],c[28]);
//50 - 13 e
counter154 u135(p[639],p[670],p[701],p[732],p[763],p[794],p[825],p[856],p[887],p[918],p[949],p[980],p[1011],o3[32],o2[33],o0[35],o1[35],o2[35],o3[35]);
ha u136(Cout[34],o1[34],s[29],c[29]);
//51 - 12 e
counter53 u137(p[671],p[702],p[733],p[764],p[795],s1[35],c1[35],Cout[35]);
counter53 u138(p[826],p[857],p[888],p[919],p[950],s1[36],c1[36],Cout[36]);
counter53 u139(p[981],p[1012],o3[33],o2[34],o1[35],s1[37],c1[37],Cout[37]);
//52 - 11 e
counter53 u140(p[703],p[734],p[765],p[796],p[827],s1[38],c1[38],Cout[38]);
counter53 u141(p[858],p[889],p[920],p[951],p[982],s1[39],c1[39],Cout[39]);
counter53 u142(p[1013],o3[34],o2[35],c1[35],c1[36],s1[40],c1[40],Cout[40]);
//53 -10 e
counter53 u143(p[735],p[766],p[797],p[828],p[859],s1[41],c1[41],Cout[41]);
counter53 u144(p[890],p[921],p[952],p[983],p[1014],s1[42],c1[42],Cout[42]);
counter53 u145(o3[35],Cout[35],Cout[36],Cout[37],c1[38],s1[43],c1[43],Cout[43]);
//54- 9 e
counter53 u146(p[767],p[798],p[829],p[860],p[891],s1[44],c1[44],Cout[44]);
counter53 u147(p[922],p[953],p[984],p[1015],Cout[38],s1[45],c1[45],Cout[45]);
fa u148(Cout[39],Cout[40],c1[41],s[30],c[30]);
//55 - 8 e
counter53 u149(p[799],p[830],p[861],p[892],p[923],s1[46],c1[46],Cout[46]);
counter53 u150(p[954],p[985],p[1016],Cout[41],Cout[42],s1[47],c1[47],Cout[47]);
fa u151(Cout[43],c1[44],c1[45],s[31],c[31]);
//56 - 7 e
counter53 u152(p[831],p[862],p[893],p[924],p[955],s1[48],c1[48],Cout[48]);
counter53 u153(p[986],p[1017],Cout[44],Cout[45],c1[46],s1[49],c1[49],Cout[49]);
ha u154(c1[47],c[31],s[32],c[32]);
//57 - 6 e
counter53 u155(p[863],p[894],p[925],p[956],p[987],s1[50],c1[50],Cout[50]);
counter53 u156(p[1018],Cout[46],Cout[47],c1[48],c1[49],s1[51],c1[51],Cout[51]);
//56 - 5 e
counter53 u157(p[895],p[926],p[957],p[988],p[1019],s1[52],c1[52],Cout[52]);
fa u158(Cout[48],Cout[49],c1[50],s[33],c[33]);
//57 - 4 e
counter53 u159(p[927],p[958],p[989],p[1020],Cout[50],s1[53],c1[53],Cout[53]);
fa u160(Cout[51],c1[52],c[33],s[34],c[34]);
//58 - 3 e
counter53 u161(p[959],p[990],p[1021],Cout[52],c1[53],s1[54],c1[54],Cout[54]);
//59 - 2e
fa u162(p[991],p[1022],Cout[53],s[35],c[35]);
//62 - 1 e
fa u163(p[1023],Cout[54],c[35],s[36],c[36]);

//second stage
//0
ha u164(p[0],c[36],s[37],c[37]);
//1//
fa u165(p[1],p[32],c[37],s[38],c[38]);
//2//
fa u166(p[2],p[33],c[38],s[39],c[39]);
//3//
fa u167(p[3],p[34],p[65],s[40],c[40]);
//4
fa u168(s[12],p[66],p[97],s[41],c[41]);
//5
ha u169(s1[0],p[129],s[42],c[42]);
//6
counter53 u170(s1[1],p[130],p[161],p[192],c[42],s1[55],c1[55],Cout[55]);
//7
counter53 u171(s1[2],s[13],p[193],p[224],c1[55],s1[56],c1[56],Cout[56]);
//8
counter53 u172(s1[3],s1[4],p[225],p[256],Cout[55],s1[57],c1[57],Cout[57]);
//9
counter53 u173(s1[5],s1[6],p[226],p[257],Cout[56],s1[58],c1[58],Cout[58]);
//10
counter53 u174(s1[7],s1[8],s[14],p[258],Cout[57],s1[59],c1[59],Cout[59]);
ha u175(p[289],c1[58],s[43],c[43]);
//11
counter53 u176(s1[9],s1[10],s[15],p[259],Cout[58],s1[60],c1[60],Cout[60]);
fa u177(p[290],p[321],c1[59],s[44],c[44]);
//12
counter53 u178(o0[0],c1[9],c1[10],c[15],Cout[59],s1[61],c1[61],Cout[61]);
//13
fa u179(o0[1],Cout[9],Cout[10],s[45],c[45]);
//14
fa u180(o0[2],o2[0],o1[1],s[46],c[46]);
//15
fa u181(o0[3],s[16],o2[1],s[47],c[47]);
//16
counter53 u182(o0[4],s[17],o2[2],o1[3],c[47],s1[62],c1[62],Cout[62]);
//17
counter53 u183(o0[5],s[18],o3[2],o2[3],c1[62],s1[63],c1[63],Cout[63]);
//18
counter53 u184(o0[6],s1[11],o2[4],o1[5],Cout[62],s1[64],c1[64],Cout[64]);
//19
counter53 u185(o0[7],s1[12],o3[4],o2[5],Cout[63],s1[65],c1[65],Cout[65]);
//20
counter53 u186(o0[8],s1[13],s[19],Cout[11],Cout[64],s1[66],c1[66],Cout[66]);
//21
counter53 u187(o0[9],s1[14],s[20],o2[7],Cout[12],s1[67],c1[67],Cout[67]);
counter53 u188(o1[8],c1[13],c[19],Cout[65],c1[66],s1[68],c1[68],Cout[68]);
//22
counter53 u189(o0[10],s1[15],s[21],o3[7],o2[8],s1[69],c1[69],Cout[69]);
counter53 u190(Cout[13],o1[9],c1[14],c[20],Cout[66],s1[70],c1[70],Cout[70]);
ha u191(c1[67],c1[68],s[48],c[48]);
//23
counter154 u192(o0[11],s1[16],s[22],p[736],o3[8],o2[9],Cout[14],o1[10],c1[15],c[21],Cout[67],Cout[68],c1[69],c1[70],c[48],o0[36],o1[36],o2[36],o3[36]);
//24
counter53 u193(o0[12],s1[17],s[23],p[737],p[768],s1[71],c1[71],Cout[71]);
counter53 u194(o3[9],o2[10],Cout[15],o1[11],c1[16],s1[72],c1[72],Cout[72]);
fa u195(c[22],Cout[69],Cout[70],s[49],c[49]);
//25
counter154 u196(o0[13],s1[18],s[24],p[738],p[769],p[800],o3[10],o2[11],Cout[16],o1[12],c1[17],c[23],o2[36],c1[71],c1[72],o0[37],o1[37],o2[37],o3[37]);
//26
counter154 u197(o0[14],s1[19],s[25],p[739],p[770],p[801],p[832],o3[11],o2[12],Cout[17],o1[13],c1[18],c[24],o3[36],Cout[71],o0[38],o1[38],o2[38],o3[38]);
//27
fa u198(O0[0],s[26],c[25],s[50],c[50]);
//28
ha u199(O0[1],o3[37],s[51],c[51]);
//29
ha u200(O0[2],O1[1],s[52],c[52]);
//30
fa u201(O0[3],O3[0],O2[1],s[53],c[53]);
//31
counter53 u202(O0[4],p[992],O4[0],O3[1],O2[2],s1[73],c1[73],Cout[73]);
//32
counter53 u203(O0[5],O4[1],O3[2],O2[3],c1[73],s1[74],c1[74],Cout[74]);
//33
counter53 u204(O0[6],O3[3],O2[4],O1[5],Cout[73],s1[75],c1[75],Cout[75]);
//34
counter53 u205(O0[7],O2[5],O1[6],Cout[74],c1[75],s1[76],c1[76],Cout[76]);
//35
counter53 u206(o0[15],o0[16],O2[6],O1[7],Cout[75],s1[77],c1[77],Cout[77]);
//36
counter53 u207(o0[17],o0[18],o1[15],o1[16],Cout[76],s1[78],c1[78],Cout[78]);
//37
counter53 u208(o0[19],o0[20],o1[17],o1[18],Cout[77],s1[79],c1[79],Cout[79]);
//38
counter53 u209(o0[21],o0[22],o1[19],o1[20],Cout[78],s1[80],c1[80],Cout[80]);
//39
fa u210(o0[23],o0[24],Cout[79],s[54],c[54]);
//40
counter53 u211(o0[25],s1[20],s1[21],o2[21],o2[22],s1[81],c1[81],Cout[81]);
fa u212(o1[23],o1[24],Cout[80],s[55],c[55]);
//41
counter53 u213(o0[26],s1[22],s1[23],o2[24],o1[25],s1[82],c1[82],Cout[82]);
fa u214(c1[20],c1[21],c1[81],s[56],c[56]);
//42
counter53 u215(o0[27],s1[24],s1[25],Cout[21],o1[26],s1[83],c1[83],Cout[83]);
counter53 u216(c1[22],c1[23],Cout[81],c1[82],c[56],s1[84],c1[84],Cout[84]);
//43
counter53 u217(o0[28],s1[26],s1[27],c1[24],c1[25],s1[85],c1[85],Cout[85]);
fa u218(Cout[82],c1[83],c1[84],s[57],c[57]);
//44
counter53 u219(o0[29],s1[28],s1[29],c1[27],Cout[83],s1[86],c1[86],Cout[86]);
fa u220(Cout[84],c1[85],c[57],s[58],c[58]);
//45
counter53 u221(o0[30],s1[30],s1[31],Cout[85],c1[86],s1[87],c1[87],Cout[87]);
//46
counter53 u222(o0[31],s1[32],s[26],c1[31],Cout[86],s1[88],c1[88],Cout[88]);
//47
counter53 u223(o0[32],s1[33],s[27],c[26],Cout[87],s1[89],c1[89],Cout[89]);
//48
counter53 u224(o0[33],s1[34],c[27],Cout[88],c1[89],s1[90],c1[90],Cout[90]);
//49
counter53 u225(o0[34],s[28],c1[34],Cout[89],c1[90],s1[91],c1[91],Cout[91]);
//50
counter53 u226(o0[35],s[29],c[28],Cout[90],c1[91],s1[92],c1[92],Cout[92]);
//51
counter53 u227(s1[35],s1[36],s1[37],c[29],Cout[91],s1[93],c1[93],Cout[93]);
//52
counter53 u228(s1[38],s1[39],s1[40],c1[37],Cout[92],s1[94],c1[94],Cout[94]);
//53
counter53 u229(s1[41],s1[42],s1[43],c1[39],c1[40],s1[95],c1[95],Cout[95]);
ha u230(Cout[93],c1[94],s[59],c[59]);
//54
counter53 u231(s1[44],s1[45],s[30],c1[42],c1[43],s1[96],c1[96],Cout[96]);
fa u232(Cout[94],c1[95],c[59],s[60],c[60]);
//55
counter53 u233(s1[46],s1[47],s[31],c[30],Cout[95],s1[97],c1[97],Cout[97]);
ha u234(c1[96],c[60],s[61],c[61]);
//56
counter53 u235(s1[48],s1[49],s[32],Cout[96],c1[97],s1[98],c1[98],Cout[98]);
//57
counter53 u236(s1[50],s1[51],c[32],Cout[97],c1[98],s1[99],c1[99],Cout[99]);
//58
counter53 u237(s1[52],s[33],c1[51],Cout[98],c1[99],s1[100],c1[100],Cout[100]);
//59
fa u238(s1[53],s[34],Cout[99],s[62],c[62]);
//60
fa u239(s1[54],c[34],Cout[100],s[63],c[63]);
//61
fa u240(s[35],c1[54],c[63],s[64],c[64]);
//62
ha u241(s[36],c[64],s[65],c[65]);

//third stage
//0
ha u242(s[37],c[65],s[66],c[66]);
//1
ha u243(s[38],c[66],s[67],c[67]);
//2
fa u244(s[39],p[64],c[67],s[68],c[68]);
//3
fa u245(s[40],c[39],p[96],s[69],c[69]);
//4
fa u246(s[41],c[40],p[128],s[70],c[70]);
//5
fa u247(s[42],c[41],p[160],s[71],c[71]);
//6
ha u248(s1[55],c[71],s[72],c[72]);
//7
ha u249(s1[56],c[72],s[73],c[73]);
//8
fa u250(s1[57],c1[56],c[73],s[74],c[74]);
//9
fa u251(s1[58],c1[57],p[288],s[75],c[75]);
//10
fa u252(s1[59],s[43],p[320],s[76],c[76]);
//11
counter53 u253(s1[60],s[44],p[352],c[43],c[76],s1[101],c1[101],Cout[101]);
//12
fa u254(s1[61],c1[60],c[44],s[77],c[77]);
//13
counter53 u255(s[45],c1[61],Cout[60],Cout[101],c[77],s1[102],c1[102],Cout[102]);
//14
fa u256(s[46],Cout[61],c[45],s[78],c[78]);
//15
counter53 u257(s[47],c[46],o3[0],Cout[102],c[78],s1[103],c1[103],Cout[103]);
//16
fa u258(s1[62],c[16],c1[103],s[79],c[79]);
//17
counter53 u259(s1[63],o1[4],c[17],Cout[103],c[79],s1[104],c1[104],Cout[104]);
//18
fa u260(s1[64],c1[63],c[18],s[80],c[80]);
//19
counter53 u261(s1[65],c1[64],o1[6],c1[11],Cout[104],s1[105],c1[105],Cout[105]);
//20
counter53 u262(s1[66],c1[65],o1[7],c1[12],c1[105],s1[106],c1[106],Cout[106]);
//21
fa u263(s1[67],s1[68],Cout[105],s[81],c[81]);
//22
counter53 u264(s1[69],s1[70],s[48],Cout[106],c[81],s1[107],c1[107],Cout[107]);
//23
ha u265(o0[36],c1[107],s[82],c[82]);
//24
counter53 u266(s1[71],s1[72],s[49],o1[36],Cout[107],s1[108],c1[108],Cout[108]);
//25
fa u267(o0[37],c[49],c1[108],s[83],c[83]);
//26
counter53 u268(o0[38],Cout[72],o1[37],Cout[108],c[83],s1[109],c1[109],Cout[109]);
//27
fa u269(s[50],o2[37],o1[38],s[84],c[84]);
//28
counter53 u270(s[51],o2[38],c[50],Cout[109],c[84],s1[110],c1[110],Cout[110]);
//29
fa u271(s[52],o3[38],c[51],s[85],c[85]);
//30
counter53 u272(s[53],c[52],O1[2],Cout[110],c[85],s1[111],c1[111],Cout[111]);
//31
fa u273(s1[73],c[53],O1[3],s[86],c[86]);
//32
fa u274(s1[74],O1[4],Cout[111],s[87],c[87]);
//33
fa u275(s1[75],c1[74],c[87],s[88],c[88]);
//34
ha u276(s1[76],c[88],s[89],c[89]);
//35
fa u277(s1[77],c1[76],c[89],s[90],c[90]);
//36
fa u278(s1[78],c1[77],c[90],s[91],c[91]);
//37
fa u279(s1[79],c1[78],c[91],s[92],c[92]);
//38
fa u280(s1[80],c1[79],c[92],s[93],c[93]);
//39
fa u281(s[54],c1[80],c[93],s[94],c[94]);
//40
fa u282(s1[81],s[55],c[54],s[95],c[95]);
//41
fa u283(s1[82],s[56],c[55],s[96],c[96]);
//42
fa u284(s1[83],s1[84],c[96],s[97],c[97]);
//43
fa u285(s1[85],s[57],c[97],s[98],c[98]);
//44
fa u286(s1[86],s[58],c[98],s[99],c[99]);
//45
fa u287(s1[87],c[58],c[99],s[100],c[100]);
//46
fa u288(s1[88],c1[87],c[100],s[101],c[101]);
//47
fa u289(s1[89],c1[88],c[101],s[102],c[102]);
//48
ha u290(s1[90],c[102],s[103],c[103]);
//49
ha u291(s1[91],c[103],s[104],c[104]);
//50
ha u292(s1[92],c[104],s[105],c[105]);
//51
fa u293(s1[93],c1[92],c[105],s[106],c[106]);
//52
fa u294(s1[94],c1[93],c[106],s[107],c[107]);
//53
fa u295(s1[95],s[59],c[107],s[108],c[108]);
//54
fa u296(s1[96],s[60],c[108],s[109],c[109]);
//55
fa u297(s1[97],s[61],c[109],s[110],c[110]);
//56
fa u298(s1[98],c[61],c[110],s[111],c[111]);
//57
ha u299(s1[99],c[111],s[112],c[112]);
//58
ha u300(s1[100],c[112],s[113],c[113]);
//59
fa u301(s[62],c1[100],c[113],s[114],c[114]);
//60
fa u302(s[63],c[62],c[114],s[115],c[115]);
//61
ha u303(s[64],c[115],s[116],c[116]);
//62
ha u304(s[65],c[116],s[117],c[117]);

//final stage
//0
ha u305(s[66],c[117],y[0],c[118]);
//1
ha u306(s[67],c[118],y[1],c[119]);
//2
ha u307(s[68],c[119],y[2],c[120]);
//3
fa u308(s[69],c[68],c[120],y[3],c[121]);
//4
fa u309(s[70],c[69],c[121],y[4],c[122]);
//5
fa u310(s[71],c[70],c[122],y[5],c[123]);
//6
ha u311(s[72],c[123],y[6],c[124]);
//7
ha u312(s[73],c[124],y[7],c[125]);
//8
ha u313(s[74],c[125],y[8],c[126]);
//9
fa u314(s[75],c[74],c[126],y[9],c[127]);
//10
fa u315(s[76],c[75],c[127],y[10],c[128]);
//11
ha u316(s1[101],c[128],y[11],c[129]);
//12
fa u317(s[77],c1[101],c[129],y[12],c[130]);
//13
ha u318(s1[102],c[130],y[13],c[131]);
//14
fa u319(s[78],c1[102],c[131],y[14],c[132]);
//15
ha u320(s1[103],c[132],y[15],c[133]);
//16
ha u321(s[79],c[133],y[16],c[134]);
//17
ha u322(s1[104],c[134],y[17],c[135]);
//18
fa u323(s[80],c1[104],c[135],y[18],c[136]);
//19
fa u324(s1[105],c[80],c[136],y[19],c[137]);
//20
ha u325(s1[106],c[137],y[20],c[138]);
//21
fa u326(s[81],c1[106],c[138],y[21],c[139]);
//22
ha u327(s1[107],c[139],y[22],c[140]);
//23
ha u328(s[82],c[140],y[23],c[141]);
//24
fa u329(s1[108],c[82],c[141],y[24],c[142]);
//25
ha u330(s[83],c[142],y[25],c[143]);
//26
ha u331(s1[109],c[143],y[26],c[144]);
//27
fa u332(s[84],c1[109],c[144],y[27],c[145]);
//28
ha u333(s1[110],c[145],y[28],c[146]);
//29
fa u334(s[85],c1[110],c[146],y[29],c[147]);
//30
ha u335(s1[111],c[147],y[30],c[148]);
//31
fa u336(s[86],c1[111],c[148],y[31],c[149]);
//32
fa u337(s[87],c[86],c[149],y[32],c[150]);
//33
ha u338(s[88],c[150],y[33],c[151]);
//34
ha u339(s[89],c[151],y[34],c[152]);
//35
ha u340(s[90],c[152],y[35],c[153]);
//36
ha u341(s[91],c[153],y[36],c[154]);
//37
ha u342(s[92],c[154],y[37],c[155]);
//38
ha u343(s[93],c[155],y[38],c[156]);
//39
ha u344(s[94],c[156],y[39],c[157]);
//40
fa u345(s[95],c[94],c[157],y[40],c[158]);
//41
fa u346(s[96],c[95],c[158],y[41],c[159]);
//42
ha u347(s[97],c[159],y[42],c[160]);
//43
ha u348(s[98],c[160],y[43],c[161]);
//44
ha u349(s[99],c[161],y[44],c[162]);
//45
ha u350(s[100],c[162],y[45],c[163]);
//46
ha u351(s[101],c[163],y[46],c[164]);
//47
ha u352(s[102],c[164],y[47],c[165]);
//48
ha u353(s[103],c[165],y[48],c[166]);
//49
ha u354(s[104],c[166],y[49],c[167]);
//50
ha u355(s[105],c[167],y[50],c[168]);
//51
ha u356(s[106],c[168],y[51],c[169]);
//52
ha u357(s[107],c[169],y[52],c[170]);
//53
ha u358(s[108],c[170],y[53],c[171]);
//54
ha u359(s[109],c[171],y[54],c[172]);
//55
ha u360(s[110],c[172],y[55],c[173]);
//56
ha u361(s[111],c[173],y[56],c[174]);
//57
ha u362(s[112],c[174],y[57],c[175]);
//58
ha u363(s[113],c[175],y[58],c[176]);
//59
ha u364(s[114],c[176],y[59],c[177]);
//60
ha u365(s[115],c[177],y[60],c[178]);
//61
ha u366(s[116],c[178],y[61],c[179]);
//62
ha u367(s[117],c[179],y[62],c[180]);

        
assign c[180] = y[63];

endmodule

module counter315(i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,O0,O1,O2,O3,O4);
input i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30;
  output O0,O1,O2,O3,O4;
  wire s[11:8];
  wire c[11:8];
  wire o0[1:0],o1[1:0],o2[1:0],o3[1:0];
 
  counter154 u11(i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,o0[0],o1[0],o2[0],o3[0]);
  counter154 u12(i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,o0[1],o1[1],o2[1],o3[1]);
 
fa u13(i30,o0[1],o0[0],s[8],c[8]);
fa u14(o1[0],o1[1],c[8],s[9],c[9]);
fa u15(o2[0],o2[1],c[9],s[10],c[10]);
fa u16(o3[0],o3[1],c[10],s[11],c[11]);
 
  assign s[8]=O0;
  assign s[9]=O1;
  assign s[10]=O2;
  assign s[11]=O3;
  assign c[11]=O4;
endmodule
  
module counter154(Z0,Z1,Z2,Z3,Z4,Z5,Z6,Z7,Z8,Z9,Z10,Z11,Z12,Z13,Z14,o0,o1,o2,o3);
input Z0,Z1,Z2,Z3,Z4,Z5,Z6,Z7,Z8,Z9,Z10,Z11,Z12,Z13,Z14;
output o0,o1,o2,o3;
wire s[7:0];
wire c[7:0];
wire [1:0]s1,c1,Cout;


fa u1(Z0,Z1,Z2,s[0],c[0]);
fa u2(Z3,Z4,Z5,s[1],c[1]);
fa u3(Z6,Z7,Z8,s[2],c[2]);
fa u4(Z9,Z10,Z11,s[3],c[3]);
fa u5(Z12,Z13,Z14,s[4],c[4]);

counter53 u6(s[0],s[1],s[2],s[3],s[4],s1[0],c1[0],Cout[0]);
counter53 u7(c[0],c[1],c[2],c[3],c[4],s1[1],c1[1],Cout[1]);

assign s1[0]=o0;
ha u8(c1[0],s1[1],s[5],c[5]);
fa u9(Cout[0],c1[1],c[0],s[6],c[6]);
ha u10(Cout[1],c[1],s[7],c[7]);
assign s[5] = o1;
assign s[6] = o2;
assign s[7] = o3;
endmodule  

module counter53(X0,X1,X2,X3,X4,s1,c1,Cout);
input X0,X1,X2,X3,X4;
output s1,c1,Cout;
wire Y[4:0],P,R;
wire R1,R2,P1,P2;
wire t1,t2,t3;

assign Y[0] = X3 | X4;
assign Y[1] = X3 & X4;
assign Y[2] = X1 | X2;
assign Y[3] = X1 & X2;
assign Y[4] = X0;
assign R1 = Y[0] & ~Y[1];
assign R2 = Y[2] & ~Y[3];
assign R = R1 ^ R2 ;
assign P1 = ~R & Y[3];
assign P2 = R & Y[4];
assign P = P1 | P2;
assign t1 = Y[1] | Y[2];
assign t2 = Y[0] & t1;
assign Cout = t2 & P;
assign t3 = Y[0] & t1;
assign c1 = t3 ^ P; 
assign s1 = R ^ Y[4];

endmodule

module fa(a,b,c,s,co);
input a,b,c;
output s,co;
assign s = a ^ b ^ c;
assign co = (a & b) | (b & c) | (c & a);
endmodule

module ha(a,b,s,c);
input a,b;
output s,c;
assign s = a ^ b;
assign c = a & b;
endmodule 

module mul_16x16(a,b,p);
input [15:0]a,b;
output [255:0]p;

mul_8x8 u31(a[7:0],b[7:0],p[63:0]);
mul_8x8 u32(a[15:8],b[7:0],p[127:64]);
mul_8x8 u33(a[7:0],b[15:8],p[191:128]);
mul_8x8 u34(a[15:8],b[15:8],p[255:192]);

endmodule

module mul_8x8(a,b,p);
input [7:0]a,b;
output [63:0]p;

mul_4x4 u27(a[3:0],b[3:0],p[15:0]);
mul_4x4 u28(a[7:4],b[3:0],p[31:16]);
mul_4x4 u29(a[3:0],b[7:4],p[47:32]);
mul_4x4 u30(a[7:4],b[7:4],p[63:48]);

endmodule


module mul_4x4(a,b,p);
input [3:0]a,b;
output [15:0]p;

and u11(p[0],a[0],b[0]);
and u12(p[1],a[1],b[0]);
and u13(p[2],a[2],b[0]);
and u14(p[3],a[3],b[0]);
and u15(p[4],a[0],b[1]);
and u16(p[5],a[1],b[1]);
and u17(p[6],a[2],b[1]);
and u18(p[7],a[3],b[1]);
and u19(p[8],a[0],b[2]);
and u20(p[9],a[1],b[2]);
and u21(p[10],a[2],b[2]);
and u22(p[11],a[3],b[2]);
and u23(p[12],a[0],b[3]);
and u24(p[13],a[1],b[3]);
and u25(p[14],a[2],b[3]);
and u26(p[15],a[3],b[3]);

endmodule

`default_nettype wire
